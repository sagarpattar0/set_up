sagar.sv
