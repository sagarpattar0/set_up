hd bsjdjbnisdsad
